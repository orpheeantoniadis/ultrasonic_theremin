// nios.v

// Generated using ACDS version 17.0 595

`timescale 1 ps / 1 ps
module nios (
		input  wire        clk_clk,                    //               clk.clk
		output wire        i2s0_export_mck,            //       i2s0_export.mck
		output wire        i2s0_export_lrck,           //                  .lrck
		output wire        i2s0_export_data,           //                  .data
		output wire        i2s0_export_sck,            //                  .sck
		output wire [7:0]  led_sel_b_export_readdata,  //  led_sel_b_export.readdata
		output wire [7:0]  led_sel_g_export_readdata,  //  led_sel_g_export.readdata
		output wire [7:0]  led_sel_r_export_readdata,  //  led_sel_r_export.readdata
		output wire [11:0] led_selc_n_export_readdata, // led_selc_n_export.readdata
		output wire [7:0]  ledsa_export_export,        //      ledsa_export.export
		output wire [7:0]  ledsb_export_export,        //      ledsb_export.export
		input  wire        reset_reset_n,              //             reset.reset_n
		input  wire        ultrasound_export_echo,     // ultrasound_export.echo
		output wire        ultrasound_export_trig      //                  .trig
	);

	wire         altpll_0_c0_clk;                                           // altpll_0:c0 -> [I2S_0:clock, mm_interconnect_0:altpll_0_c0_clk, rst_controller:clk]
	wire  [31:0] cpu_data_master_readdata;                                  // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire         cpu_data_master_waitrequest;                               // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire         cpu_data_master_debugaccess;                               // cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire  [15:0] cpu_data_master_address;                                   // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                                // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire         cpu_data_master_read;                                      // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire         cpu_data_master_readdatavalid;                             // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire         cpu_data_master_write;                                     // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire  [31:0] cpu_data_master_writedata;                                 // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                           // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire         cpu_instruction_master_waitrequest;                        // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire  [15:0] cpu_instruction_master_address;                            // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire         cpu_instruction_master_read;                               // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire         cpu_instruction_master_readdatavalid;                      // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;    // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest; // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire         mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire         mm_interconnect_0_ultrasound_0_avalon_slave_0_chipselect;  // mm_interconnect_0:ultrasound_0_avalon_slave_0_chipselect -> ultrasound_0:ChipSelect
	wire  [31:0] mm_interconnect_0_ultrasound_0_avalon_slave_0_readdata;    // ultrasound_0:ReadData -> mm_interconnect_0:ultrasound_0_avalon_slave_0_readdata
	wire         mm_interconnect_0_ultrasound_0_avalon_slave_0_read;        // mm_interconnect_0:ultrasound_0_avalon_slave_0_read -> ultrasound_0:Read
	wire         mm_interconnect_0_ledmatrix_0_avalon_slave_0_chipselect;   // mm_interconnect_0:ledmatrix_0_avalon_slave_0_chipselect -> ledmatrix_0:ChipSelect
	wire  [15:0] mm_interconnect_0_ledmatrix_0_avalon_slave_0_readdata;     // ledmatrix_0:ReadData -> mm_interconnect_0:ledmatrix_0_avalon_slave_0_readdata
	wire   [6:0] mm_interconnect_0_ledmatrix_0_avalon_slave_0_address;      // mm_interconnect_0:ledmatrix_0_avalon_slave_0_address -> ledmatrix_0:Address
	wire         mm_interconnect_0_ledmatrix_0_avalon_slave_0_read;         // mm_interconnect_0:ledmatrix_0_avalon_slave_0_read -> ledmatrix_0:Read
	wire         mm_interconnect_0_ledmatrix_0_avalon_slave_0_write;        // mm_interconnect_0:ledmatrix_0_avalon_slave_0_write -> ledmatrix_0:Write
	wire  [15:0] mm_interconnect_0_ledmatrix_0_avalon_slave_0_writedata;    // mm_interconnect_0:ledmatrix_0_avalon_slave_0_writedata -> ledmatrix_0:WriteData
	wire         mm_interconnect_0_i2s_0_avalon_slave_0_chipselect;         // mm_interconnect_0:I2S_0_avalon_slave_0_chipselect -> I2S_0:chip_select
	wire   [2:0] mm_interconnect_0_i2s_0_avalon_slave_0_address;            // mm_interconnect_0:I2S_0_avalon_slave_0_address -> I2S_0:addresse
	wire         mm_interconnect_0_i2s_0_avalon_slave_0_write;              // mm_interconnect_0:I2S_0_avalon_slave_0_write -> I2S_0:write
	wire  [15:0] mm_interconnect_0_i2s_0_avalon_slave_0_writedata;          // mm_interconnect_0:I2S_0_avalon_slave_0_writedata -> I2S_0:write_data
	wire  [31:0] mm_interconnect_0_sys_id_control_slave_readdata;           // Sys_ID:readdata -> mm_interconnect_0:Sys_ID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sys_id_control_slave_address;            // mm_interconnect_0:Sys_ID_control_slave_address -> Sys_ID:address
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;            // cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;         // cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;         // mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;             // mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;                // mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;          // mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;               // mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;           // mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_readdata;             // altpll_0:readdata -> mm_interconnect_0:altpll_0_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_altpll_0_pll_slave_address;              // mm_interconnect_0:altpll_0_pll_slave_address -> altpll_0:address
	wire         mm_interconnect_0_altpll_0_pll_slave_read;                 // mm_interconnect_0:altpll_0_pll_slave_read -> altpll_0:read
	wire         mm_interconnect_0_altpll_0_pll_slave_write;                // mm_interconnect_0:altpll_0_pll_slave_write -> altpll_0:write
	wire  [31:0] mm_interconnect_0_altpll_0_pll_slave_writedata;            // mm_interconnect_0:altpll_0_pll_slave_writedata -> altpll_0:writedata
	wire         mm_interconnect_0_onchip_ram_s1_chipselect;                // mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_readdata;                  // onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	wire  [11:0] mm_interconnect_0_onchip_ram_s1_address;                   // mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	wire   [3:0] mm_interconnect_0_onchip_ram_s1_byteenable;                // mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	wire         mm_interconnect_0_onchip_ram_s1_write;                     // mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	wire  [31:0] mm_interconnect_0_onchip_ram_s1_writedata;                 // mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	wire         mm_interconnect_0_onchip_ram_s1_clken;                     // mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	wire         mm_interconnect_0_ledsa_s1_chipselect;                     // mm_interconnect_0:ledsA_s1_chipselect -> ledsA:chipselect
	wire  [31:0] mm_interconnect_0_ledsa_s1_readdata;                       // ledsA:readdata -> mm_interconnect_0:ledsA_s1_readdata
	wire   [1:0] mm_interconnect_0_ledsa_s1_address;                        // mm_interconnect_0:ledsA_s1_address -> ledsA:address
	wire         mm_interconnect_0_ledsa_s1_write;                          // mm_interconnect_0:ledsA_s1_write -> ledsA:write_n
	wire  [31:0] mm_interconnect_0_ledsa_s1_writedata;                      // mm_interconnect_0:ledsA_s1_writedata -> ledsA:writedata
	wire         mm_interconnect_0_timer_0_s1_chipselect;                   // mm_interconnect_0:timer_0_s1_chipselect -> timer_0:chipselect
	wire  [15:0] mm_interconnect_0_timer_0_s1_readdata;                     // timer_0:readdata -> mm_interconnect_0:timer_0_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_0_s1_address;                      // mm_interconnect_0:timer_0_s1_address -> timer_0:address
	wire         mm_interconnect_0_timer_0_s1_write;                        // mm_interconnect_0:timer_0_s1_write -> timer_0:write_n
	wire  [15:0] mm_interconnect_0_timer_0_s1_writedata;                    // mm_interconnect_0:timer_0_s1_writedata -> timer_0:writedata
	wire         mm_interconnect_0_ledsb_s1_chipselect;                     // mm_interconnect_0:ledsB_s1_chipselect -> ledsB:chipselect
	wire  [31:0] mm_interconnect_0_ledsb_s1_readdata;                       // ledsB:readdata -> mm_interconnect_0:ledsB_s1_readdata
	wire   [1:0] mm_interconnect_0_ledsb_s1_address;                        // mm_interconnect_0:ledsB_s1_address -> ledsB:address
	wire         mm_interconnect_0_ledsb_s1_write;                          // mm_interconnect_0:ledsB_s1_write -> ledsB:write_n
	wire  [31:0] mm_interconnect_0_ledsb_s1_writedata;                      // mm_interconnect_0:ledsB_s1_writedata -> ledsB:writedata
	wire         irq_mapper_receiver0_irq;                                  // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                                  // timer_0:irq -> irq_mapper:receiver1_irq
	wire  [31:0] cpu_irq_irq;                                               // irq_mapper:sender_irq -> cpu:irq
	wire         rst_controller_reset_out_reset;                            // rst_controller:reset_out -> [I2S_0:nReset, mm_interconnect_0:I2S_0_reset_sink_reset_bridge_in_reset_reset]
	wire         cpu_debug_reset_request_reset;                             // cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                        // rst_controller_001:reset_out -> [Sys_ID:reset_n, altpll_0:reset, cpu:reset_n, irq_mapper:reset, jtag_uart:rst_n, ledmatrix_0:nReset, ledsA:reset_n, ledsB:reset_n, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_translator:in_reset, ultrasound_0:nReset]
	wire         rst_controller_001_reset_out_reset_req;                    // rst_controller_001:reset_req -> [cpu:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	wire         rst_controller_002_reset_out_reset;                        // rst_controller_002:reset_out -> [mm_interconnect_0:timer_0_reset_reset_bridge_in_reset_reset, timer_0:reset_n]

	i2s_controller i2s_0 (
		.addresse    (mm_interconnect_0_i2s_0_avalon_slave_0_address),    // avalon_slave_0.address
		.chip_select (mm_interconnect_0_i2s_0_avalon_slave_0_chipselect), //               .chipselect
		.write       (mm_interconnect_0_i2s_0_avalon_slave_0_write),      //               .write
		.write_data  (mm_interconnect_0_i2s_0_avalon_slave_0_writedata),  //               .writedata
		.clock       (altpll_0_c0_clk),                                   //     clock_sink.clk
		.GPIO_2_D0   (i2s0_export_mck),                                   //    conduit_end.mck
		.GPIO_2_D1   (i2s0_export_lrck),                                  //               .lrck
		.GPIO_2_D2   (i2s0_export_data),                                  //               .data
		.GPIO_2_D3   (i2s0_export_sck),                                   //               .sck
		.nReset      (~rst_controller_reset_out_reset)                    //     reset_sink.reset_n
	);

	nios_Sys_ID sys_id (
		.clock    (clk_clk),                                         //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),             //         reset.reset_n
		.readdata (mm_interconnect_0_sys_id_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sys_id_control_slave_address)   //              .address
	);

	nios_altpll_0 altpll_0 (
		.clk                (clk_clk),                                        //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),             // inclk_interface_reset.reset
		.read               (mm_interconnect_0_altpll_0_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_altpll_0_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_altpll_0_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_altpll_0_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_altpll_0_pll_slave_writedata), //                      .writedata
		.c0                 (altpll_0_c0_clk),                                //                    c0.clk
		.scandone           (),                                               //           (terminated)
		.scandataout        (),                                               //           (terminated)
		.areset             (1'b0),                                           //           (terminated)
		.locked             (),                                               //           (terminated)
		.phasedone          (),                                               //           (terminated)
		.phasecounterselect (4'b0000),                                        //           (terminated)
		.phaseupdown        (1'b0),                                           //           (terminated)
		.phasestep          (1'b0),                                           //           (terminated)
		.scanclk            (1'b0),                                           //           (terminated)
		.scanclkena         (1'b0),                                           //           (terminated)
		.scandata           (1'b0),                                           //           (terminated)
		.configupdate       (1'b0)                                            //           (terminated)
	);

	nios_cpu cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.d_readdatavalid                     (cpu_data_master_readdatavalid),                     //                          .readdatavalid
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.i_readdatavalid                     (cpu_instruction_master_readdatavalid),              //                          .readdatavalid
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	nios_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                   //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	LedMatrix #(
		.size (16)
	) ledmatrix_0 (
		.Clk        (clk_clk),                                                 //          clock.clk
		.Address    (mm_interconnect_0_ledmatrix_0_avalon_slave_0_address),    // avalon_slave_0.address
		.ChipSelect (mm_interconnect_0_ledmatrix_0_avalon_slave_0_chipselect), //               .chipselect
		.Read       (mm_interconnect_0_ledmatrix_0_avalon_slave_0_read),       //               .read
		.Write      (mm_interconnect_0_ledmatrix_0_avalon_slave_0_write),      //               .write
		.ReadData   (mm_interconnect_0_ledmatrix_0_avalon_slave_0_readdata),   //               .readdata
		.WriteData  (mm_interconnect_0_ledmatrix_0_avalon_slave_0_writedata),  //               .writedata
		.nReset     (~rst_controller_001_reset_out_reset),                     //     reset_sink.reset_n
		.LED_SelC_n (led_selc_n_export_readdata),                              //     LED_SelC_n.readdata
		.LED_Sel_B  (led_sel_b_export_readdata),                               //      LED_Sel_B.readdata
		.LED_Sel_G  (led_sel_g_export_readdata),                               //      LED_Sel_G.readdata
		.LED_Sel_R  (led_sel_r_export_readdata)                                //      LED_Sel_R.readdata
	);

	nios_ledsA ledsa (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_ledsa_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledsa_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledsa_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledsa_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledsa_s1_readdata),   //                    .readdata
		.out_port   (ledsa_export_export)                    // external_connection.export
	);

	nios_ledsA ledsb (
		.clk        (clk_clk),                               //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),   //               reset.reset_n
		.address    (mm_interconnect_0_ledsb_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_ledsb_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_ledsb_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_ledsb_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_ledsb_s1_readdata),   //                    .readdata
		.out_port   (ledsb_export_export)                    // external_connection.export
	);

	nios_onchip_ram onchip_ram (
		.clk        (clk_clk),                                    //   clk1.clk
		.address    (mm_interconnect_0_onchip_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),         // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req),     //       .reset_req
		.freeze     (1'b0)                                        // (terminated)
	);

	nios_timer_0 timer_0 (
		.clk        (clk_clk),                                 //   clk.clk
		.reset_n    (~rst_controller_002_reset_out_reset),     // reset.reset_n
		.address    (mm_interconnect_0_timer_0_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_0_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_0_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_0_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_0_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver1_irq)                 //   irq.irq
	);

	Ultrasound ultrasound_0 (
		.Clk        (clk_clk),                                                  //          clock.clk
		.ChipSelect (mm_interconnect_0_ultrasound_0_avalon_slave_0_chipselect), // avalon_slave_0.chipselect
		.Read       (mm_interconnect_0_ultrasound_0_avalon_slave_0_read),       //               .read
		.ReadData   (mm_interconnect_0_ultrasound_0_avalon_slave_0_readdata),   //               .readdata
		.nReset     (~rst_controller_001_reset_out_reset),                      //     reset_sink.reset_n
		.Echo       (ultrasound_export_echo),                                   //    conduit_end.echo
		.Trig       (ultrasound_export_trig)                                    //               .trig
	);

	nios_mm_interconnect_0 mm_interconnect_0 (
		.altpll_0_c0_clk                              (altpll_0_c0_clk),                                           //                            altpll_0_c0.clk
		.clk_0_clk_clk                                (clk_clk),                                                   //                              clk_0_clk.clk
		.cpu_reset_reset_bridge_in_reset_reset        (rst_controller_001_reset_out_reset),                        //        cpu_reset_reset_bridge_in_reset.reset
		.I2S_0_reset_sink_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                            // I2S_0_reset_sink_reset_bridge_in_reset.reset
		.timer_0_reset_reset_bridge_in_reset_reset    (rst_controller_002_reset_out_reset),                        //    timer_0_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                      (cpu_data_master_address),                                   //                        cpu_data_master.address
		.cpu_data_master_waitrequest                  (cpu_data_master_waitrequest),                               //                                       .waitrequest
		.cpu_data_master_byteenable                   (cpu_data_master_byteenable),                                //                                       .byteenable
		.cpu_data_master_read                         (cpu_data_master_read),                                      //                                       .read
		.cpu_data_master_readdata                     (cpu_data_master_readdata),                                  //                                       .readdata
		.cpu_data_master_readdatavalid                (cpu_data_master_readdatavalid),                             //                                       .readdatavalid
		.cpu_data_master_write                        (cpu_data_master_write),                                     //                                       .write
		.cpu_data_master_writedata                    (cpu_data_master_writedata),                                 //                                       .writedata
		.cpu_data_master_debugaccess                  (cpu_data_master_debugaccess),                               //                                       .debugaccess
		.cpu_instruction_master_address               (cpu_instruction_master_address),                            //                 cpu_instruction_master.address
		.cpu_instruction_master_waitrequest           (cpu_instruction_master_waitrequest),                        //                                       .waitrequest
		.cpu_instruction_master_read                  (cpu_instruction_master_read),                               //                                       .read
		.cpu_instruction_master_readdata              (cpu_instruction_master_readdata),                           //                                       .readdata
		.cpu_instruction_master_readdatavalid         (cpu_instruction_master_readdatavalid),                      //                                       .readdatavalid
		.altpll_0_pll_slave_address                   (mm_interconnect_0_altpll_0_pll_slave_address),              //                     altpll_0_pll_slave.address
		.altpll_0_pll_slave_write                     (mm_interconnect_0_altpll_0_pll_slave_write),                //                                       .write
		.altpll_0_pll_slave_read                      (mm_interconnect_0_altpll_0_pll_slave_read),                 //                                       .read
		.altpll_0_pll_slave_readdata                  (mm_interconnect_0_altpll_0_pll_slave_readdata),             //                                       .readdata
		.altpll_0_pll_slave_writedata                 (mm_interconnect_0_altpll_0_pll_slave_writedata),            //                                       .writedata
		.cpu_debug_mem_slave_address                  (mm_interconnect_0_cpu_debug_mem_slave_address),             //                    cpu_debug_mem_slave.address
		.cpu_debug_mem_slave_write                    (mm_interconnect_0_cpu_debug_mem_slave_write),               //                                       .write
		.cpu_debug_mem_slave_read                     (mm_interconnect_0_cpu_debug_mem_slave_read),                //                                       .read
		.cpu_debug_mem_slave_readdata                 (mm_interconnect_0_cpu_debug_mem_slave_readdata),            //                                       .readdata
		.cpu_debug_mem_slave_writedata                (mm_interconnect_0_cpu_debug_mem_slave_writedata),           //                                       .writedata
		.cpu_debug_mem_slave_byteenable               (mm_interconnect_0_cpu_debug_mem_slave_byteenable),          //                                       .byteenable
		.cpu_debug_mem_slave_waitrequest              (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),         //                                       .waitrequest
		.cpu_debug_mem_slave_debugaccess              (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),         //                                       .debugaccess
		.I2S_0_avalon_slave_0_address                 (mm_interconnect_0_i2s_0_avalon_slave_0_address),            //                   I2S_0_avalon_slave_0.address
		.I2S_0_avalon_slave_0_write                   (mm_interconnect_0_i2s_0_avalon_slave_0_write),              //                                       .write
		.I2S_0_avalon_slave_0_writedata               (mm_interconnect_0_i2s_0_avalon_slave_0_writedata),          //                                       .writedata
		.I2S_0_avalon_slave_0_chipselect              (mm_interconnect_0_i2s_0_avalon_slave_0_chipselect),         //                                       .chipselect
		.jtag_uart_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //            jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),       //                                       .write
		.jtag_uart_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),        //                                       .read
		.jtag_uart_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                                       .readdata
		.jtag_uart_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                                       .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                                       .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  //                                       .chipselect
		.ledmatrix_0_avalon_slave_0_address           (mm_interconnect_0_ledmatrix_0_avalon_slave_0_address),      //             ledmatrix_0_avalon_slave_0.address
		.ledmatrix_0_avalon_slave_0_write             (mm_interconnect_0_ledmatrix_0_avalon_slave_0_write),        //                                       .write
		.ledmatrix_0_avalon_slave_0_read              (mm_interconnect_0_ledmatrix_0_avalon_slave_0_read),         //                                       .read
		.ledmatrix_0_avalon_slave_0_readdata          (mm_interconnect_0_ledmatrix_0_avalon_slave_0_readdata),     //                                       .readdata
		.ledmatrix_0_avalon_slave_0_writedata         (mm_interconnect_0_ledmatrix_0_avalon_slave_0_writedata),    //                                       .writedata
		.ledmatrix_0_avalon_slave_0_chipselect        (mm_interconnect_0_ledmatrix_0_avalon_slave_0_chipselect),   //                                       .chipselect
		.ledsA_s1_address                             (mm_interconnect_0_ledsa_s1_address),                        //                               ledsA_s1.address
		.ledsA_s1_write                               (mm_interconnect_0_ledsa_s1_write),                          //                                       .write
		.ledsA_s1_readdata                            (mm_interconnect_0_ledsa_s1_readdata),                       //                                       .readdata
		.ledsA_s1_writedata                           (mm_interconnect_0_ledsa_s1_writedata),                      //                                       .writedata
		.ledsA_s1_chipselect                          (mm_interconnect_0_ledsa_s1_chipselect),                     //                                       .chipselect
		.ledsB_s1_address                             (mm_interconnect_0_ledsb_s1_address),                        //                               ledsB_s1.address
		.ledsB_s1_write                               (mm_interconnect_0_ledsb_s1_write),                          //                                       .write
		.ledsB_s1_readdata                            (mm_interconnect_0_ledsb_s1_readdata),                       //                                       .readdata
		.ledsB_s1_writedata                           (mm_interconnect_0_ledsb_s1_writedata),                      //                                       .writedata
		.ledsB_s1_chipselect                          (mm_interconnect_0_ledsb_s1_chipselect),                     //                                       .chipselect
		.onchip_ram_s1_address                        (mm_interconnect_0_onchip_ram_s1_address),                   //                          onchip_ram_s1.address
		.onchip_ram_s1_write                          (mm_interconnect_0_onchip_ram_s1_write),                     //                                       .write
		.onchip_ram_s1_readdata                       (mm_interconnect_0_onchip_ram_s1_readdata),                  //                                       .readdata
		.onchip_ram_s1_writedata                      (mm_interconnect_0_onchip_ram_s1_writedata),                 //                                       .writedata
		.onchip_ram_s1_byteenable                     (mm_interconnect_0_onchip_ram_s1_byteenable),                //                                       .byteenable
		.onchip_ram_s1_chipselect                     (mm_interconnect_0_onchip_ram_s1_chipselect),                //                                       .chipselect
		.onchip_ram_s1_clken                          (mm_interconnect_0_onchip_ram_s1_clken),                     //                                       .clken
		.Sys_ID_control_slave_address                 (mm_interconnect_0_sys_id_control_slave_address),            //                   Sys_ID_control_slave.address
		.Sys_ID_control_slave_readdata                (mm_interconnect_0_sys_id_control_slave_readdata),           //                                       .readdata
		.timer_0_s1_address                           (mm_interconnect_0_timer_0_s1_address),                      //                             timer_0_s1.address
		.timer_0_s1_write                             (mm_interconnect_0_timer_0_s1_write),                        //                                       .write
		.timer_0_s1_readdata                          (mm_interconnect_0_timer_0_s1_readdata),                     //                                       .readdata
		.timer_0_s1_writedata                         (mm_interconnect_0_timer_0_s1_writedata),                    //                                       .writedata
		.timer_0_s1_chipselect                        (mm_interconnect_0_timer_0_s1_chipselect),                   //                                       .chipselect
		.ultrasound_0_avalon_slave_0_read             (mm_interconnect_0_ultrasound_0_avalon_slave_0_read),        //            ultrasound_0_avalon_slave_0.read
		.ultrasound_0_avalon_slave_0_readdata         (mm_interconnect_0_ultrasound_0_avalon_slave_0_readdata),    //                                       .readdata
		.ultrasound_0_avalon_slave_0_chipselect       (mm_interconnect_0_ultrasound_0_avalon_slave_0_chipselect)   //                                       .chipselect
	);

	nios_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),  // reset_in1.reset
		.clk            (altpll_0_c0_clk),                //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),          // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
